/*
E/16/070
DE SILVA N.S.C.K.S.
LAB05 PART2_TESTBENCH
*/

// testbench for register file
module reg_file_tb;
    
    reg [7:0] WRITEDATA;
    reg [2:0] WRITEREG, READREG1, READREG2;
    reg CLK, RESET, WRITEENABLE; 
    wire [7:0] REGOUT1, REGOUT2;
    
    reg_file myregfile(WRITEDATA, REGOUT1, REGOUT2, WRITEREG, READREG1, READREG2, WRITEENABLE, CLK, RESET);
       
    initial
    begin
        CLK = 1'b1;
        
        // generate files needed to plot the waveform using GTKWave
        $dumpfile("reg_file_wavedata.vcd");
		$dumpvars(0, reg_file_tb);
        
        // assign values with time to input signals to see output 
        RESET = 1'b0;
        WRITEENABLE = 1'b0;
        
        #1
        RESET = 1'b1;
        READREG1 = 3'd2;
        READREG2 = 3'd6;
        
        #8
        RESET = 1'b0;
        
        #5
        WRITEREG = 3'd7;
        WRITEDATA = 8'd17;
        WRITEENABLE = 1'b1;
        
        #10
        WRITEENABLE = 1'b0;
        
        #2
        READREG1 = 3'd7;
        
        #9
        WRITEREG = 3'd2;
        WRITEDATA = 8'd37;
        WRITEENABLE = 1'b1;
        READREG1 = 3'd2;
	RESET = 1'b1 ;

	#10
	RESET = 1'b0 ;
        
        #6
        WRITEENABLE = 1'b1;

        #6
        WRITEREG = 3'd6;
        WRITEDATA = 8'd47;
        WRITEENABLE = 1'b1;
        READREG2 = 3'd6;
        
        #10
        WRITEDATA = 8'd97;
        WRITEENABLE = 1'b1;
        READREG2 = 3'd6;
        
        #10
        WRITEENABLE = 1'b0;
        
        #6
        WRITEREG = 3'd5;
        WRITEDATA = 8'd57;
        WRITEENABLE = 1'b1;
        
        #5
        WRITEENABLE = 1'b0;
        
        #2
        WRITEREG = 3'd3;
        WRITEDATA = 8'd45;
        WRITEENABLE = 1'b1;
        READREG2 = 3'd3;	
	
	#10
        $finish;
    end
    
    // clock signal generation
    always
        #5 CLK = ~CLK;
        

endmodule
